// ECE423_QSYS_sram.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module ECE423_QSYS_sram (
		output wire [0:0]  bridge_memory_tcm_chipselect_n_out,   // bridge.memory_tcm_chipselect_n_out
		output wire [1:0]  bridge_memory_tcm_byteenable_n_out,   //       .memory_tcm_byteenable_n_out
		output wire [18:0] bridge_memory_tcm_address_out,        //       .memory_tcm_address_out
		inout  wire [15:0] bridge_memory_tcm_data_out,           //       .memory_tcm_data_out
		output wire [0:0]  bridge_memory_tcm_write_n_out,        //       .memory_tcm_write_n_out
		output wire [0:0]  bridge_memory_tcm_outputenable_n_out, //       .memory_tcm_outputenable_n_out
		input  wire        clk_clk,                              //    clk.clk
		input  wire        reset_reset_n,                        //  reset.reset_n
		input  wire [18:0] uas_address,                          //    uas.address
		input  wire [1:0]  uas_burstcount,                       //       .burstcount
		input  wire        uas_read,                             //       .read
		input  wire        uas_write,                            //       .write
		output wire        uas_waitrequest,                      //       .waitrequest
		output wire        uas_readdatavalid,                    //       .readdatavalid
		input  wire [1:0]  uas_byteenable,                       //       .byteenable
		output wire [15:0] uas_readdata,                         //       .readdata
		input  wire [15:0] uas_writedata,                        //       .writedata
		input  wire        uas_lock,                             //       .lock
		input  wire        uas_debugaccess                       //       .debugaccess
	);

	wire         memory_sharer_tcm_request;                           // memory_sharer:request -> memory_bridge:request
	wire  [15:0] memory_sharer_tcm_memory_tcm_data_out_out;           // memory_sharer:memory_tcm_data_out -> memory_bridge:tcs_memory_tcm_data_out
	wire   [0:0] memory_sharer_tcm_memory_tcm_write_n_out_out;        // memory_sharer:memory_tcm_write_n_out -> memory_bridge:tcs_memory_tcm_write_n_out
	wire  [15:0] memory_sharer_tcm_memory_tcm_data_out_in;            // memory_bridge:tcs_memory_tcm_data_in -> memory_sharer:memory_tcm_data_in
	wire         memory_sharer_tcm_memory_tcm_data_out_outen;         // memory_sharer:memory_tcm_data_outen -> memory_bridge:tcs_memory_tcm_data_outen
	wire   [0:0] memory_sharer_tcm_memory_tcm_chipselect_n_out_out;   // memory_sharer:memory_tcm_chipselect_n_out -> memory_bridge:tcs_memory_tcm_chipselect_n_out
	wire         memory_sharer_tcm_grant;                             // memory_bridge:grant -> memory_sharer:grant
	wire   [0:0] memory_sharer_tcm_memory_tcm_outputenable_n_out_out; // memory_sharer:memory_tcm_outputenable_n_out -> memory_bridge:tcs_memory_tcm_outputenable_n_out
	wire  [18:0] memory_sharer_tcm_memory_tcm_address_out_out;        // memory_sharer:memory_tcm_address_out -> memory_bridge:tcs_memory_tcm_address_out
	wire   [1:0] memory_sharer_tcm_memory_tcm_byteenable_n_out_out;   // memory_sharer:memory_tcm_byteenable_n_out -> memory_bridge:tcs_memory_tcm_byteenable_n_out
	wire         memory_tcm_data_outen;                               // memory:tcm_data_outen -> memory_sharer:tcs0_data_outen
	wire         memory_tcm_outputenable_n_out;                       // memory:tcm_outputenable_n_out -> memory_sharer:tcs0_outputenable_n_out
	wire         memory_tcm_request;                                  // memory:tcm_request -> memory_sharer:tcs0_request
	wire   [1:0] memory_tcm_byteenable_n_out;                         // memory:tcm_byteenable_n_out -> memory_sharer:tcs0_byteenable_n_out
	wire         memory_tcm_write_n_out;                              // memory:tcm_write_n_out -> memory_sharer:tcs0_write_n_out
	wire         memory_tcm_grant;                                    // memory_sharer:tcs0_grant -> memory:tcm_grant
	wire         memory_tcm_chipselect_n_out;                         // memory:tcm_chipselect_n_out -> memory_sharer:tcs0_chipselect_n_out
	wire  [18:0] memory_tcm_address_out;                              // memory:tcm_address_out -> memory_sharer:tcs0_address_out
	wire  [15:0] memory_tcm_data_out;                                 // memory:tcm_data_out -> memory_sharer:tcs0_data_out
	wire  [15:0] memory_tcm_data_in;                                  // memory_sharer:tcs0_data_in -> memory:tcm_data_in
	wire         rst_controller_reset_out_reset;                      // rst_controller:reset_out -> [memory:reset_reset, memory_bridge:reset, memory_sharer:reset_reset]

	ECE423_QSYS_sram_memory #(
		.TCM_ADDRESS_W                  (19),
		.TCM_DATA_W                     (16),
		.TCM_BYTEENABLE_W               (2),
		.TCM_READ_WAIT                  (10),
		.TCM_WRITE_WAIT                 (10),
		.TCM_SETUP_WAIT                 (10),
		.TCM_DATA_HOLD                  (10),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (2),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (0),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (1),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (1),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (0),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (1),
		.ACTIVE_LOW_OUTPUTENABLE        (1),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) memory (
		.clk_clk                (clk_clk),                        //   clk.clk
		.reset_reset            (rst_controller_reset_out_reset), // reset.reset
		.uas_address            (uas_address),                    //   uas.address
		.uas_burstcount         (uas_burstcount),                 //      .burstcount
		.uas_read               (uas_read),                       //      .read
		.uas_write              (uas_write),                      //      .write
		.uas_waitrequest        (uas_waitrequest),                //      .waitrequest
		.uas_readdatavalid      (uas_readdatavalid),              //      .readdatavalid
		.uas_byteenable         (uas_byteenable),                 //      .byteenable
		.uas_readdata           (uas_readdata),                   //      .readdata
		.uas_writedata          (uas_writedata),                  //      .writedata
		.uas_lock               (uas_lock),                       //      .lock
		.uas_debugaccess        (uas_debugaccess),                //      .debugaccess
		.tcm_write_n_out        (memory_tcm_write_n_out),         //   tcm.write_n_out
		.tcm_chipselect_n_out   (memory_tcm_chipselect_n_out),    //      .chipselect_n_out
		.tcm_outputenable_n_out (memory_tcm_outputenable_n_out),  //      .outputenable_n_out
		.tcm_request            (memory_tcm_request),             //      .request
		.tcm_grant              (memory_tcm_grant),               //      .grant
		.tcm_address_out        (memory_tcm_address_out),         //      .address_out
		.tcm_byteenable_n_out   (memory_tcm_byteenable_n_out),    //      .byteenable_n_out
		.tcm_data_out           (memory_tcm_data_out),            //      .data_out
		.tcm_data_outen         (memory_tcm_data_outen),          //      .data_outen
		.tcm_data_in            (memory_tcm_data_in)              //      .data_in
	);

	ECE423_QSYS_sram_memory_bridge memory_bridge (
		.clk                               (clk_clk),                                             //   clk.clk
		.reset                             (rst_controller_reset_out_reset),                      // reset.reset
		.request                           (memory_sharer_tcm_request),                           //   tcs.request
		.grant                             (memory_sharer_tcm_grant),                             //      .grant
		.tcs_memory_tcm_chipselect_n_out   (memory_sharer_tcm_memory_tcm_chipselect_n_out_out),   //      .memory_tcm_chipselect_n_out_out
		.tcs_memory_tcm_byteenable_n_out   (memory_sharer_tcm_memory_tcm_byteenable_n_out_out),   //      .memory_tcm_byteenable_n_out_out
		.tcs_memory_tcm_address_out        (memory_sharer_tcm_memory_tcm_address_out_out),        //      .memory_tcm_address_out_out
		.tcs_memory_tcm_data_out           (memory_sharer_tcm_memory_tcm_data_out_out),           //      .memory_tcm_data_out_out
		.tcs_memory_tcm_data_outen         (memory_sharer_tcm_memory_tcm_data_out_outen),         //      .memory_tcm_data_out_outen
		.tcs_memory_tcm_data_in            (memory_sharer_tcm_memory_tcm_data_out_in),            //      .memory_tcm_data_out_in
		.tcs_memory_tcm_write_n_out        (memory_sharer_tcm_memory_tcm_write_n_out_out),        //      .memory_tcm_write_n_out_out
		.tcs_memory_tcm_outputenable_n_out (memory_sharer_tcm_memory_tcm_outputenable_n_out_out), //      .memory_tcm_outputenable_n_out_out
		.memory_tcm_chipselect_n_out       (bridge_memory_tcm_chipselect_n_out),                  //   out.memory_tcm_chipselect_n_out
		.memory_tcm_byteenable_n_out       (bridge_memory_tcm_byteenable_n_out),                  //      .memory_tcm_byteenable_n_out
		.memory_tcm_address_out            (bridge_memory_tcm_address_out),                       //      .memory_tcm_address_out
		.memory_tcm_data_out               (bridge_memory_tcm_data_out),                          //      .memory_tcm_data_out
		.memory_tcm_write_n_out            (bridge_memory_tcm_write_n_out),                       //      .memory_tcm_write_n_out
		.memory_tcm_outputenable_n_out     (bridge_memory_tcm_outputenable_n_out)                 //      .memory_tcm_outputenable_n_out
	);

	ECE423_QSYS_sram_memory_sharer memory_sharer (
		.clk_clk                       (clk_clk),                                             //   clk.clk
		.reset_reset                   (rst_controller_reset_out_reset),                      // reset.reset
		.request                       (memory_sharer_tcm_request),                           //   tcm.request
		.grant                         (memory_sharer_tcm_grant),                             //      .grant
		.memory_tcm_address_out        (memory_sharer_tcm_memory_tcm_address_out_out),        //      .memory_tcm_address_out_out
		.memory_tcm_byteenable_n_out   (memory_sharer_tcm_memory_tcm_byteenable_n_out_out),   //      .memory_tcm_byteenable_n_out_out
		.memory_tcm_outputenable_n_out (memory_sharer_tcm_memory_tcm_outputenable_n_out_out), //      .memory_tcm_outputenable_n_out_out
		.memory_tcm_write_n_out        (memory_sharer_tcm_memory_tcm_write_n_out_out),        //      .memory_tcm_write_n_out_out
		.memory_tcm_data_out           (memory_sharer_tcm_memory_tcm_data_out_out),           //      .memory_tcm_data_out_out
		.memory_tcm_data_in            (memory_sharer_tcm_memory_tcm_data_out_in),            //      .memory_tcm_data_out_in
		.memory_tcm_data_outen         (memory_sharer_tcm_memory_tcm_data_out_outen),         //      .memory_tcm_data_out_outen
		.memory_tcm_chipselect_n_out   (memory_sharer_tcm_memory_tcm_chipselect_n_out_out),   //      .memory_tcm_chipselect_n_out_out
		.tcs0_request                  (memory_tcm_request),                                  //  tcs0.request
		.tcs0_grant                    (memory_tcm_grant),                                    //      .grant
		.tcs0_address_out              (memory_tcm_address_out),                              //      .address_out
		.tcs0_byteenable_n_out         (memory_tcm_byteenable_n_out),                         //      .byteenable_n_out
		.tcs0_outputenable_n_out       (memory_tcm_outputenable_n_out),                       //      .outputenable_n_out
		.tcs0_write_n_out              (memory_tcm_write_n_out),                              //      .write_n_out
		.tcs0_data_out                 (memory_tcm_data_out),                                 //      .data_out
		.tcs0_data_in                  (memory_tcm_data_in),                                  //      .data_in
		.tcs0_data_outen               (memory_tcm_data_outen),                               //      .data_outen
		.tcs0_chipselect_n_out         (memory_tcm_chipselect_n_out)                          //      .chipselect_n_out
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
